`timescale 1ns/10ps

`include "UART_TX_2.v"

module UART_TB ();

  // Testbench uses a 25 MHz clock
  // Want to interface to 115200 baud UART
  // 25000000 / 115200 = 217 Clocks Per Bit.
  parameter c_CLOCK_PERIOD_NS = 40;
  parameter c_CLKS_PER_BIT    = 217;
  parameter c_BIT_PERIOD      = 8600;
  
  reg r_Clock = 0;
  reg clk_in = 0;
  reg r_TX_DV = 0;
  wire w_TX_Active, w_UART_Line;
  wire w_TX_Serial;
  reg [7:0] r_TX_Byte = 0;
  wire [7:0] w_RX_Byte;

  UART_RX #(.cpb(c_CLKS_PER_BIT)) UART_RX_Inst
    (.clk(r_Clock),
     .rx_data_in(w_UART_Line),
     .rx_dv(w_RX_DV),
     .rx_data_out(w_RX_Byte)
     );
  
  UART_TX #(.cpb(c_CLKS_PER_BIT)) UART_TX_Inst
    (.clk(r_Clock),
     .tx_dv(r_TX_DV),
     .tx_data_in(r_TX_Byte),
     .tx_active(w_TX_Active),
     .tx_data_out(w_TX_Serial),
     .tx_done()
     );
	BRG B1 (.clk_in(clk_in), .clk_out(r_clk));

  // Keeps the UART Receive input high (default) when
  // UART transmitter is not active
  assign w_UART_Line = w_TX_Active ? w_TX_Serial : 1'b1;
    
  always
    #(c_CLOCK_PERIOD_NS/2) r_Clock <= !r_Clock;
  
  // Main Testing:
  initial
    begin
      // Tell UART to send a command (exercise TX)
      //@(posedge r_Clock); 
      
      @(posedge r_Clock);
	begin
     	r_TX_DV   <= 1'b1;
 	r_TX_Byte <= 8'h69;
     	
	end
	 @(posedge r_Clock);
     	begin
	r_TX_DV <= 1'b0;
	end
	 
      // Check that the correct command was received
      @(posedge w_RX_DV);
	begin
	
      if (w_RX_Byte == 8'h69)
        $display($time,"Test Passed - Correct Byte Received");
      else
        $display("Test Failed - Incorrect Byte Received");
	end
      $finish();
    end
endmodule

